module roi_axis(
  
  input logic xy_0_i,
  input logic xy_1_i


);
  
endmodule