module roi_apb(
  input logic xy_0_o,
  input logic xy_1_o
);
  
endmodule