module roi_apb(
  input   logic         clk_i,
  input   logic         arst_i,

  

  output  logic  [31:0] xy_0_o,
  output  logic  [31:0] xy_1_o
);
  
endmodule