`timescale 1ns / 1ps

module roi_top_tb();





endmodule
