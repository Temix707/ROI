`timescale 1ns / 1ps

module roi_axis_tb();





endmodule
