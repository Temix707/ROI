`timescale 1ns / 1ps

module roi_apb_tb();





endmodule
